-- revision history:
-- 06.07.2015     Alex Schönberger    created


entity tb_alu is
end entity tb_alu;

architecture behav_tb_alu of tb_alu is

  component alu 
  end component alu;

  --signal 

begin

--  uut: alu
--    PORT MAP(
--    );

  process
  begin

    wait;
  end process;

end architecture behav_tb_alu;
