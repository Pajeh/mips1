library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library WORK;
use WORK.cpu_pack.all;

entity tb_fsm2 is
end entity tb_fsm2;

architecture behavioural of tb_fsm2 is
end architecture;