-- revision history:
-- 06.07.2015     Alex Schönberger    created

entity cpu_datapath is

end entity cpu_datapath;


architecture structure_cpu_datapath of cpu_datapath is

begin

end architecture structure_cpu_datapath;