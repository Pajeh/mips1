-- revision history:
-- 03.08.2015     Patrick Appenheimer    created

entity tb_execution is
end entity tb_execution;

architecture behav_tb_execution of tb_execution is
begin

end architecture behav_tb_execution;
