-- revision history:
-- 06.07.2015     Alex Schönberger    created

entity cpu_control is

end entity cpu_control;


architecture structure_cpu_control of cpu_control is

begin

end architecture structure_cpu_control;